module gameController (clk, reset, enable, gameLevel, userWon, signalLess, signalGreater, userPrimeNbrTensDgt, userPrimeNbrUnitsDgt);
	input clk, reset, enable;
	input [3:0] userPrimeNbrTensDgt, userPrimeNbrUnitsDgt;	
	input [1:0] gameLevel;
	output userWon, signalLess, signalGreater;

	wire [6:0] randomPrimeNbr;
	reg [6:0] userPrimeNbr;

	LFSR_Prime inst_RndmPrimeGenerator (
		.clk (clk)
		, .rst (reset)
		, .gameLevel (gameLevel)
		, .enable (enable)
		, .Q_out (randomPrimeNbr)
	);

	always @ (posedge clk)
	begin
		if (userPrimeNbrTensDgt >= 10 && userPrimeNbrUnitsDgt >= 10 )
		begin
			userPrimeNbr <= 99;
		end
		else if (userPrimeNbrTensDgt >= 10 )
		begin
			userPrimeNbr <= 90 + userPrimeNbrUnitsDgt;
		end
		else if (userPrimeNbrUnitsDgt >= 10 )
		begin
			userPrimeNbr <= userPrimeNbrTensDgt + 9;
		end
		else 
		begin
			userPrimeNbr <= 10*userPrimeNbrTensDgt + userPrimeNbrUnitsDgt;
		end
	end

	always @ (posedge clk)
	begin
		if (reset == 1'b0)
		begin
			signalLess <= 1'b0;
			signalGreater <= 1'b0;
			userWon <= 1'b0;
		end
		else
		begin
			// logic to compare the random prime number with the
			// generated prime number.
			if (randomPrimeNbr == userPrimeNbr)
			begin
				userWon <= 1'b1;
			end
			// check to see if the random number that the user
			// input is less than the one generated by the FPGA,
			// if yes, then turn on the 'signalLess' LED.
			else if (randomPrimeNbr < userPrimeNbr)
			begin
				signalLess <= 1'b1;
			end
			// check to see if the random number from the user is
			// greater than the prime number generated. If yes,
			// then turn on the 'signalGreater' LED.
			else if (randomPrimeNbr > userPrimeNbr)
			begin
				signalGreater <= 1'b1;
			end
		end
	end
endmodule
	
