module checkPassword(clk,rst,Load_Button_PSWD_Game_Control,Logout_Pulse,Data_in,Authenticated,Logout_RED, access_allowed, userUniqueID);
	input clk,rst;
	input Load_Button_PSWD_Game_Control,Logout_Pulse; // Load_Button_PSWD_Game_Control ouput pulse from the button shaper
	input [3:0]Data_in; // data enetered using the switches
//	input [15:0] ROM_Password; // input from the Multi_Password_ROM
	reg [2:0] ROM_Address; // output to Multi_Password_ROM
	output reg Authenticated,Logout_RED, access_allowed; // Authentication
	
	wire [15:0] ROM_PeopleSoftID, ROM_Password;
	reg [3:0] STATE;
	reg [15:0] Password_Entered;
	output reg [2:0] userUniqueID;
	reg peopleSoftIDStage;
	
	parameter [3:0]
		Digit1 = 0,Digit2 = 1,Digit3 = 2,Digit4 = 3,
		Fetch_ROM_Data = 4, Wait1 = 5, Wait2 = 6,ROM_DATA_READ = 7, CheckPassword = 8,
		Authorize = 9,Initial = 10, Logout_State = 11;
	
	
	always @ (posedge clk)
	begin
			access_allowed <= Authenticated;
	end
	
	// instantiate the 1-port ROM to read the user ID that the user
	// inputs.
	multiID instMultipleID (
		.address (ROM_Address),
		.clock (clk),
		.q (ROM_PeopleSoftID)
	);
	
	// Instantiate the 1-port ROM to read the password associated with
	// selected user Profile
	multiPSWD instUsrPswd (
		.address (ROM_Address),
		.clock (clk),
		.q (ROM_Password)
	);
	
	
	
	always @(posedge clk) begin
		// reset stage
			if (rst == 1'b0) begin
				Authenticated <= 1'b0;
				STATE <= Initial;
				ROM_Address <= 3'b000;
				Logout_RED <=1'b1;
				Password_Entered <= 0;
				userUniqueID <= 3'b000;
				peopleSoftIDStage <= 1'b0;
			end
			
			else begin
				case (STATE)
	// initial conditions
				Initial: begin
							peopleSoftIDStage <= 1'b0;
							userUniqueID <= 3'b000;
							Authenticated <= 1'b0;
							Logout_RED <= 1'b1;
							ROM_Address <= 3'b000;
							STATE <= Digit1;
				end
	// storing the msb bit 15-12 in Password_Entered buffer		
				Digit1: begin
							if (Load_Button_PSWD_Game_Control == 1'b1) begin
								Password_Entered[15:12] <= Data_in;
								STATE <= Digit2;
							end
							else begin
								STATE <= Digit1;
							end	
				end	
	//storing the bit from 11-8 in Password_Entered buffer
				Digit2: begin
							if (Load_Button_PSWD_Game_Control == 1'b1) begin
								Password_Entered[11:8] <= Data_in;
								STATE <= Digit3;
							end
							else begin
								STATE <= Digit2;
							end	
				end		
	// storing the bit from 7-4 in Password_Entered buffer	
				Digit3: begin
							if (Load_Button_PSWD_Game_Control == 1'b1) begin
								Password_Entered[7:4] <= Data_in;
								STATE <= Digit4;
							end
							else begin
								STATE <= Digit3;
							end	
				end	
	// storing the bit from 3-0 in Password_Entered buffer
				Digit4: begin
							if (Load_Button_PSWD_Game_Control == 1'b1) begin
								Password_Entered[3:0] <= Data_in;
								STATE <= Fetch_ROM_Data;
							end
							else begin
								STATE <= Digit4;
							end	
				end

	//first wait stage to read the data from ROM	
				
				Fetch_ROM_Data:	begin
							STATE <= Wait1;
				end
	//second wait stage			
				Wait1: begin
							STATE <= Wait2;
				end
	//third wait stage			
				Wait2: begin
						if (peopleSoftIDStage == 1'b0)
						begin
							STATE <= ROM_DATA_READ;
						end
						else begin
							STATE <= CheckPassword;
						end
				end
	// reading the data from ROM. if the password entered by the player does not match the address of the
	// ROM is incremented for 4 times and still it does not match player has to enter the correct password.
	// If the password matches it will send a signal saying that the system has been authenticated. The Authenticated
	// signal is sent to the Game_Control module.
			
				ROM_DATA_READ: begin
//						ROM_PeopleSoftID <= ROM_Password;
							
						if (Password_Entered == ROM_PeopleSoftID) begin
								userUniqueID <= ROM_Address;
								peopleSoftIDStage <= 1'b1;
								STATE <= Digit1;
						end
						else begin
							if (ROM_Address !=4) begin
								ROM_Address <= ROM_Address + 1'b1;
								STATE <= Fetch_ROM_Data;
							end
							else begin
									STATE <= Digit1;
									ROM_Address <= 3'b000;
							end
						end	
				end
				CheckPassword: begin
						if (Password_Entered == ROM_Password)
						begin
							STATE <= Authorize;
						end
						else
						begin
							STATE <= Initial;
						end
				end
				
				Authorize: begin
							Authenticated <= 1'b1;
							Logout_RED <= 1'b0;
							STATE <= Logout_State;
				end		
	// In this state the system is checking for the Logout_Pulse signal. This signal is generated by the Game 
	// acces control		
				Logout_State: begin
								if (Logout_Pulse == 0) begin
									STATE <= Logout_State;
								end
								else begin
									Authenticated <=1'b0;
									Logout_RED <= 1'b1;
									STATE <= Initial;
								end	
				end
				
				default: begin
							STATE <= Initial;
							Authenticated <= 1'b0;
							ROM_Address <= 3'b000;
							Logout_RED <= 1'b1;
				end			
				endcase
			end
		end		
endmodule
